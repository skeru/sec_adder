-- secure bit propagate generate --
library ieee;
use work.sec_type.all;
use ieee.std_logic_1164.all;

entity secure_bit_pg is
  port(
    a: in t_sec_signal;
    b: in t_sec_signal;
    rnd: in std_logic;
    p: out t_sec_signal;
    g: out t_sec_signal);
end secure_bit_pg;

architecture secure of secure_bit_pg is
  component sec_xor port(a, b: in t_sec_signal; r: in std_logic; c: out t_sec_signal); -- XOR --
  end component;
  component sec_and port(a, b: in t_sec_signal; rnd: in std_logic; c: out t_sec_signal); -- AND --
  end component;
  begin
    foo: sec_and port map (a, b, rnd, g);
    fee: sec_xor port map (a, b, rnd, p);
  end;


-- secure group propagate generate --
library ieee;
use work.sec_type.all;
use ieee.std_logic_1164.all;

entity secure_group_pg is
  port(
    p0: in t_sec_signal;
    p1: in t_sec_signal;
    g0: in t_sec_signal;
    g1: in t_sec_signal;
    rnd: in std_logic;
    p2: out t_sec_signal;
    g2: out t_sec_signal);
end secure_group_pg;

architecture secure of secure_group_pg is
  component sec_xor port(a, b: in t_sec_signal; r: in std_logic; c: out t_sec_signal); -- XOR --
  end component;
  component sec_and port(a, b: in t_sec_signal; rnd: in std_logic; c: out t_sec_signal); -- AND --
  end component;
  component sec_or port(a, b: in t_sec_signal; rnd: in std_logic; c: out t_sec_signal); -- OR --
  end component;
  signal tmp: t_sec_signal;
  begin
    foo: sec_and port map (g0, p1, rnd, tmp);
    fuu: sec_or port map (g1, tmp, rnd, g2);
    fee: sec_xor port map (p1, p0, rnd, p2);
  end;
    
-- secure group generate --
library ieee;
use work.sec_type.all;
use ieee.std_logic_1164.all;

entity secure_group_g is
  port(
    p1: in t_sec_signal;
    g0: in t_sec_signal;
    g1: in t_sec_signal;
    rnd: in std_logic;
    g2: out t_sec_signal);
end secure_group_g;

architecture secure of secure_group_g is
  component sec_and port(a, b: in t_sec_signal; rnd: in std_logic; c: out t_sec_signal); -- AND --
  end component;
  component sec_or port(a, b: in t_sec_signal; rnd: in std_logic; c: out t_sec_signal); -- OR --
  end component;
  signal tmp: t_sec_signal;
  begin
    foo: sec_and port map (g0, p1, rnd, tmp);
    fuu: sec_or port map (g1, tmp, rnd, g2);
  end;
    
-- secure Kogge Stone adder --
LIBRARY ieee;
USE ieee.std_logic_1164.all;
 
PACKAGE my_funs IS
    FUNCTION clogb2 (a: NATURAL) RETURN NATURAL;
END my_funs;
 
PACKAGE BODY my_funs IS
    FUNCTION clogb2 (a: NATURAL) RETURN NATURAL IS
        VARIABLE aggregate : NATURAL := a;
        VARIABLE return_val : NATURAL := 0;
    BEGIN
        compute_clogb2: 
        FOR i IN a DOWNTO 0 LOOP
 
            IF aggregate > 0 THEN
                return_val := return_val + 1;
            END IF;
 
            aggregate := aggregate / 2;            
        END LOOP;
 
        RETURN return_val;
 
    END clogb2;
END my_funs;
 
 
library ieee;
use ieee.std_logic_1164.all;
use work.my_funs.all;
use work.sec_type.all;

entity secure_ks_adder is
  generic( width: integer :=4);
  port(
    a: in t_sec_signal_vector(width-1 downto 0);
    b: in t_sec_signal_vector(width-1 downto 0);
    c_in: in t_sec_signal;
    rnd: in std_logic_vector(width-1 downto 0);
    sum: out t_sec_signal_vector(width-1 downto 0);
    c_out: out t_sec_signal);
end secure_ks_adder;

architecture behavioral of secure_ks_adder is
  constant depth: integer := clogb2(width);
  component sec_not port(a: in t_sec_signal; b: out t_sec_signal); -- NOT --
  end component;
  component sec_xor port(a, b: in t_sec_signal; r: in std_logic; c: out t_sec_signal); -- XOR --
  end component;
  component sec_and port(a, b: in t_sec_signal; rnd: in std_logic; c: out t_sec_signal); -- AND --
  end component;
  component secure_group_g port(p1, g0, g1: in t_sec_signal; rnd: in std_logic; g2: out t_sec_signal); -- group generate --
  end component;
  component secure_bit_pg port(a, b: in t_sec_signal; rnd: in std_logic; p, g: out t_sec_signal); -- bit generate propagate --
  end component;
  component secure_group_pg port(p0, p1, g0, g1: in t_sec_signal; rnd: in std_logic; p2, g2: out t_sec_signal); -- group generate propagate --
  end component;
  type t_adder_signal is array (depth downto 0) of t_sec_signal_vector (width-1 downto -1);
  signal p,g: t_adder_signal;
begin
  -- bit propagate and generate
  bit_propagate_generate_for: for i in width-1 downto 0 generate
    bit_map: secure_bit_pg port map (a(i), b(i), rnd(i), p(0)(i), g(0)(i));
  end generate bit_propagate_generate_for;
  p(0)(-1) <= c_in;
  g(0)(-1) <= c_in;
  --depth generation
  depth_for_gen: for d in 1 to depth generate
    constant prev: integer := d-1;
    constant shift: integer := 2**prev;
    something: for s in (-1) to d-2 generate
      p(d)(s) <= p(prev)(s);
      g(d)(s) <= g(prev)(s);      
    end generate something;
    -- group generation
    group_g_for_gen: for g_index in d-1 to (2**d)-1 generate
      group_carry_generation: secure_group_g port map (p(prev)(g_index), g(prev)(g_index-shift), g(prev)(g_index), rnd(g_index), g(d)(g_index));
    end generate group_g_for_gen;
    -- group generation and propagation
    group_gp_for_gen: for gp_index in (2**d) to width-1 generate
      group_carry_generation_propagation: secure_group_pg port map (p(prev)(gp_index-shift), p(prev)(gp_index), g(prev)(gp_index-shift), g(prev)(gp_index), rnd(gp_index), p(d)(gp_index), g(d)(gp_index));
    end generate group_gp_for_gen;
  end generate depth_for_gen;
  final_xor: for index in 0 to width-1 generate
    adder_xor: sec_xor port map (p(depth)(index), g(depth)(index-1), rnd(index), sum(index));
  end generate final_xor;
  -- carry out
  carry_out: secure_group_g port map (p(depth)(width),c_in, g(depth)(width), rnd(0), c_out);
end;